

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 2.866 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7855 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 18.299 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 88.2106 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 512.883 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2480.75 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.06379 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.356 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.71236 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.00048 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 35.013 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 168.605 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 14.176 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 68.379 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 432.958 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 2099.92 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 5.41839 LAYER VIA67 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 5.367 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8153 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 103.314 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 496.29 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA23 ;
  END SI[0]
  PIN SO[2] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 7.248 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.0553 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 55.8307 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 270.197 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 2.41472 LAYER VIA34 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 2.815 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.5402 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 103.828 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 500.616 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.07233 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.639 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.07599 LAYER METAL4 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 122.645 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 593.337 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 38.575 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 185.931 LAYER METAL5 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 565.527 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2728.02 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 2.343 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2698 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.586 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 25.688 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 123.752 LAYER METAL5 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.141 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.67821 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.969 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4733 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 1.10441 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 5.39516 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 2.114 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1683 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.844 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.682 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 24.876 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.038 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 445.159 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2158.21 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 7.45028 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 11.749 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.5127 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.1444 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.442 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.8008 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2288 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 44.6188 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 215.593 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.631119 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.663 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.0538 LAYER METAL4 ;
    ANTENNAGATEAREA 1.4638 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 50.5369 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 244.322 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.1444 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.729766 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 4.112 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1635 LAYER METAL5 ;
    ANTENNAGATEAREA 1.8317 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 85.6093 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 415.621 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.79156 LAYER VIA56 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 3.435 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5224 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1534 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 28.2876 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 132.884 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.470665 LAYER VIA23 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.729 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.50649 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.268 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48148 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 6.172 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 29.8797 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 360.281 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 1747.54 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 5.41839 LAYER VIA67 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.323 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.55363 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.55557 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2.75522 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.619 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.97739 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.55557 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2.75522 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 4.523 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7556 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 11.338 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 54.7282 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4615 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 64.7814 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 315.31 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.71384 LAYER VIA56 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.483 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9432 LAYER METAL3 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 3.991 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1967 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.188 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5267 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.586 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.41 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 132.035 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 773.314 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3733.43 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.74109 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 1.877 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.02837 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 26.836 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 129.274 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 684.421 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3305.85 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.06379 LAYER VIA56 ;
  END framing_error
END SYS_TOP

END LIBRARY
